-- a fazer
